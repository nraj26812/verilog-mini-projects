module fourbitrca (a0,b0,c0,a1,b1,a2,b2,a3,b3,s0,s111,s222,s333,c4);
input a0,b0,c0,a1,b1,a2,b2,a3,b3;
output s111,s222,s333,c4,s0;
wire s1,s2,s3,s4,s5,s6,s7,s8,s9,s10,s11,s12,c1,c2,c3;
xor(s1,a0,b0);
xor (s0,s1,c0);
and (s2,c0,s1);
and (s3,a0,b0);
or (c1,s2,c2);
xor(s4,a1,b1);
xor(s111,s4,c1);
and (s6,a1,b1);
and (s5,s4,c1);
or (c2,s5,s6);
xor(s7,a2,b2);
and (s9,a2,b2);
and (s8,s7,c2);
or (c3,s9,s8);
xor(s10,a3,b3);
xor(s222,s7,c2);
and (s11,s10, c3);
and (s12,a3,b3);
or (c4,s11,s12);
xor (s333,s10,c3);
endmodule